`ifndef __GLOBAL_CONFIG_VH__
`define __GLOBAL_CONFIG_VH__

`define PERIODS_OF_1S 50000000

`endif
